module PC_control(input C[3], input I[9], input F[3], input PC_in[16], output PC_out[16]);

endmodule;