module cpu(clk, rst_n, hlt, pc);

////////////////////////////////////////////
//IF////////////////////////////////////////
////////////////////////////////////////////



////////////////////////////////////////////
//IF/ID Reg/////////////////////////////////
////////////////////////////////////////////


////////////////////////////////////////////
//ID////////////////////////////////////////
////////////////////////////////////////////


////////////////////////////////////////////
//ID/EX Reg/////////////////////////////////
////////////////////////////////////////////


////////////////////////////////////////////
//EX////////////////////////////////////////
////////////////////////////////////////////


////////////////////////////////////////////
//EX/MEM Reg////////////////////////////////
////////////////////////////////////////////


////////////////////////////////////////////
//MEM///////////////////////////////////////
////////////////////////////////////////////


////////////////////////////////////////////
//MEM/WB Reg////////////////////////////////
////////////////////////////////////////////


////////////////////////////////////////////
//WB////////////////////////////////////////
////////////////////////////////////////////



endmodule